module or(A,B,S);
    //not and or xor 
    input A;
    input B;
    output S;

    assign S= A|B;


endmodule
