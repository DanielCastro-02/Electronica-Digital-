`timescale 1ns / 1ps
`include "sumador.v"

module sumador_tb;

	// input signals
	reg  A0;
	reg  A1;
	reg  A2;
	reg  A3;
	reg  B0;
	reg  B1;
	reg  B2;
	reg  B3;


	// output signals
	wire  S0;
	wire  S1;
	wire  S2;
	wire  S3;
	wire  Cout0;
	wire  Cout1;
	wire  Cout2;
	wire  Cout3;

// instantiation
	sumador uut(A0,B0,S0,Cout0,A1,B1,S1,Cout1,A2,B2,S2,Cout2,A3,B3,S3,Cout3);

// test vector generator
initial begin
		$dumpfile("sumador.vcd");
        $dumpvars(0,sumador_tb);
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=0;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=0;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=0;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=0;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=0;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=0;
        B2=1;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=0;
        B3=1;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=0;
        #20;
        
        A0=1;
        A1=1;
        A2=1;
        A3=1;
        B0=1;
        B1=1;
        B2=1;
        B3=1;
        #20;
        
         $display("Test complete");
end

endmodule